-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 184 04/29/2009 Service Pack 1 SJ Web Edition
-- Created on Tue Mar 16 14:21:30 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY shixu IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        tj : IN STD_LOGIC := '0';
        dp : IN STD_LOGIC := '0';
        qd : IN STD_LOGIC := '0';
        t1 : OUT STD_LOGIC;
        t2 : OUT STD_LOGIC;
        t3 : OUT STD_LOGIC;
        t4 : OUT STD_LOGIC
    );
END shixu;

ARCHITECTURE BEHAVIOR OF shixu IS
    TYPE type_fstate IS (idle,st1,s_st2,st4,st2,st3,s_st4,s_st3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,tj,dp,qd)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= idle;
            t1 <= '0';
            t2 <= '0';
            t3 <= '0';
            t4 <= '0';
        ELSE
            t1 <= '0';
            t2 <= '0';
            t3 <= '0';
            t4 <= '0';
            CASE fstate IS
                WHEN idle =>
                    IF (NOT((qd = '1'))) THEN
                        reg_fstate <= st1;
                    ELSE
                        reg_fstate <= idle;
                    END IF;

                    t1 <= '0';

                    t3 <= '0';

                    t4 <= '0';

                    t2 <= '0';
                WHEN st1 =>
                    IF (((tj = '1') AND NOT((dp = '1')))) THEN
                        reg_fstate <= st1;
                    ELSIF (((dp = '1') AND NOT((tj = '1')))) THEN
                        reg_fstate <= s_st2;
                    ELSE
                        reg_fstate <= st2;
                    END IF;

                    t1 <= '1';

                    t3 <= '0';

                    t4 <= '0';

                    t2 <= '0';
                WHEN s_st2 =>
                    IF ((tj = '1')) THEN
                        reg_fstate <= s_st2;
                    ELSE
                        reg_fstate <= s_st3;
                    END IF;

                    t1 <= '0';

                    t3 <= '0';

                    t4 <= '0';

                    t2 <= '1';
                WHEN st4 =>
                    IF (((tj = '1') AND NOT((dp = '1')))) THEN
                        reg_fstate <= st4;
                    ELSIF (((dp = '1') AND NOT((tj = '1')))) THEN
                        reg_fstate <= idle;
                    ELSE
                        reg_fstate <= st1;
                    END IF;

                    t1 <= '0';

                    t3 <= '0';

                    t4 <= '1';

                    t2 <= '0';
                WHEN st2 =>
                    IF (((tj = '1') AND NOT((dp = '1')))) THEN
                        reg_fstate <= st2;
                    ELSIF (((dp = '1') AND NOT((tj = '1')))) THEN
                        reg_fstate <= s_st3;
                    ELSE
                        reg_fstate <= st3;
                    END IF;

                    t1 <= '0';

                    t3 <= '0';

                    t4 <= '0';

                    t2 <= '1';
                WHEN st3 =>
                    IF (((tj = '1') AND NOT((dp = '1')))) THEN
                        reg_fstate <= st3;
                    ELSIF (((dp = '1') AND NOT((tj = '1')))) THEN
                        reg_fstate <= s_st4;
                    ELSE
                        reg_fstate <= st4;
                    END IF;

                    t1 <= '0';

                    t3 <= '1';

                    t4 <= '0';

                    t2 <= '0';
                WHEN s_st4 =>
                    IF ((tj = '1')) THEN
                        reg_fstate <= s_st4;
                    ELSE
                        reg_fstate <= idle;
                    END IF;

                    t1 <= '0';

                    t3 <= '0';

                    t4 <= '1';

                    t2 <= '0';
                WHEN s_st3 =>
                    IF ((tj = '1')) THEN
                        reg_fstate <= s_st3;
                    ELSE
                        reg_fstate <= s_st4;
                    END IF;

                    t1 <= '0';

                    t3 <= '1';

                    t4 <= '0';

                    t2 <= '0';
                WHEN OTHERS => 
                    t1 <= 'X';
                    t2 <= 'X';
                    t3 <= 'X';
                    t4 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
